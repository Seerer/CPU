module ALU ();
