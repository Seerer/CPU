//role as D triggers
module EX_MEM();

endmodule 